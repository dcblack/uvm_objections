`ifndef GET_ENV_SVH
`define GET_ENV_SVH
import "DPI-C" pure function string get_env(string v);
`endif
