`ifndef FORMATN_SVH
`define FORMATN_SVH
import "DPI-C" pure function string formatn(longint n);
`endif
