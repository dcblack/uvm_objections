`ifndef GET_TIME_SVH
`define GET_TIME_SVH
import "DPI-C" pure GetTimeMs64 = function longint get_time();
`endif
